module packets

pub fn hi() {
	println('hi from packets')
}